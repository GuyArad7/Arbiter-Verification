// Created by Guy Arad on 02/09/2021.

class configuration extends uvm_object;
	`uvm_object_utils(configuration)

	function new(string name = "");
		super.new(name);
	endfunction: new
endclass
