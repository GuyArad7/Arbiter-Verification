// Created by Guy Arad on 02/09/2021.

package arbiter_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "transaction.sv"
	`include "sequence_disable.sv"
	`include "sequence_read.sv"
	`include "sequence_write.sv"
	`include "sequence_random.sv"
	`include "sequence_all.sv"
	`include "sequencer.sv"
	`include "monitor_host.sv"
	`include "monitor_response.sv"
	`include "driver_host.sv"
	`include "driver_response.sv"
	`include "agent_host.sv"
	`include "agent_response.sv"
	`include "scoreboard.sv"
	`include "config.sv"
	`include "environment.sv"
	`include "test.sv"
endpackage
